module Program_Counter(
    input C_p,
    input CLK_bar,
    input CLR_bar,
    input E_p,
    output address[3:0]
    );
endmodule

module Program_Counter_tb;
endmodule
