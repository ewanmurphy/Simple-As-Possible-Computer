module Controller_Sequencer(
    input  instruction[3:0],
    output CLK,
    output CLK_bar,
    output CLR,
    output CLR_bar,
    output CON[11:0]
    );
endmodule

module Controller_Sequencer_tb;
endmodule
