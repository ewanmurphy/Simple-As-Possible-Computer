module B_Register(
    input  bus_input[7:0],
    input  L_B_bar,
    input  clk,
    output add_sub_output[7:0]
    );
endmodule

module B_Register_tb;
endmodule
