module Accumulator(bus_input, L_A_bar, E_A, CLK, bus_output, add_sub_output);
    input  [7:0] bus_input;
    input  L_A_bar;
    input  E_A;
    input  CLK;
    output [7:0] bus_output;
    output [7:0] add_sub_output;
endmodule

module Accumulator_tb;
endmodule
