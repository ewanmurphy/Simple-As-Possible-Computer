module Accumulator(
    input  bus_input[7:0],
    input  L_A_bar,
    input  E_A,
    input  clk,
    output bus_output[7:0],
    output add_sub_output[7:0]
    );
endmodule

module Accumulator_tb;
endmodule
