module Input_and_MAR(L_M_bar, CLK, bus_input, LS_output, MS_output);
    input L_M_bar;
    input CLK;
    input  [3:0] bus_input;
    output [3:0] LS_output;
    output [3:0] MS_output;
endmodule

module Input_and_MAR_tb;
endmodule
