module Output_Register(
    input L_O_bar,
    input CLK,
    input bus_input[7:0],
    output display_output[7:0]
    );
endmodule

module Output_Register_tb;
endmodule
