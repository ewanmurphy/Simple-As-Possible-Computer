module Adder_Subtractor(a_input, b_input, S_U, E_U, bus_output);
    input [7:0] a_input;
    input [7:0] b_input;
    input  S_U;
    input  E_U;
    output [7:0] bus_output;
endmodule

module Adder_Subtractor_tb;
endmodule
