module Output_Register(L_O_bar, CLK, bus_input, display_output);
    input L_O_bar;
    input CLK;
    input [7:0] bus_input;
    output [7:0] display_output;
endmodule

module Output_Register_tb;
endmodule
