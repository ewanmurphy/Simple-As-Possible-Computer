module Input_and_MAR(
    input L_M_bar,
    input CLK,
    input bus_input[3:0],
    output LS_output[3:0],
    output MS_output[3:0]
    );
endmodule

module Input_and_MAR_tb;
endmodule
