module Program_Counter(C_P, CLK_bar, CLR_bar, E_P, address);
    input C_P;
    input CLK_bar;
    input CLR_bar;
    input E_P;
    output [3:0] address;
endmodule

module Program_Counter_tb;
endmodule
