module RAM_16x8(
    input C_p,
    input CLK_bar,
    input CLR_bar,
    input E_p,
    output address[3:0]
    );
endmodule

module RAM_16x8_tb;
endmodule
