module RAM_16x8(address, data, CE_bar, memory_value);
   input [3:0] address;
   input [3:0] data;
   input CE_bar;
   output [7:0] memory_value;
endmodule

module RAM_16x8_tb;
endmodule
