module B_Register(bus_input, L_B_bar, CLK, add_sub_output);
    input [7:0] bus_input;
    input  L_B_bar;
    input  CLK;
    output [7:0] add_sub_output;
endmodule

module B_Register_tb;
endmodule
