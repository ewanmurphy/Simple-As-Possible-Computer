module Instruction_Register(
    input  L_I_bar,
    input  CLK,
    input  CLR,
    input  E_I_bar,
    input  bus_input[7:0],
    output data[3:0],
    output instruction[3:0]
    );
endmodule

module Instruction_Register_tb;
endmodule
