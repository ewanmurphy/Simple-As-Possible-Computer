module Adder_Subtractor(
    input  a_input[7:0],
    input  b_input[7:0],
    input  S_U,
    input  E_U,
    output bus_output[7:0],
    );
endmodule

module Adder_Subtractor_tb;
endmodule
